Étoile 6 br. inégales, 1 résistance

T1 1 0 2 0 Z0=120 TD=37n
T2 2 0 3 0 Z0=120 TD=41n
T3 2 0 4 0 Z0=120 TD=43n
T4 2 0 5 0 Z0=120 TD=47n
T5 2 0 6 0 Z0=120 TD=53n
T6 2 0 7 0 Z0=120 TD=59n
R2 0 3 120
VCC 1 0 PULSE(0 2 0m 1n 1n 500m)

.control
tran 10n 1000n 0 2n
plot v(6)
.endc
.end
