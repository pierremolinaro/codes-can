Ligne sans perte terminée par RC

T1 0 1 0 2 Z0=120 TD=50n
VCC 1 0 PULSE(0 5 0m 1n 1u 500m)
R1 0 2 120

.control
tran 10n 1u 0 1n
plot v(2)
.endc
.end
