Ligne sans perte ouverte

T1 0 1 0 2 Z0=120 TD=5n
VCC 1 0 PULSE(0 5 0m 1n 1n 500m)

.control
tran 10n 100n 0 1n
plot v(2)
.endc
.end
