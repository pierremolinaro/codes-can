Fermeture interrupteur sur ligne sans perte avec diodes clamping

.MODEL inter SW(RON=1m ROFF=10MEG VT=2.5 VH=.5)
.MODEL D1N4148 D (IS=0.1PA, RS=16 CJO=2PF TT=12N BV=100 IBV=0.1PA)
T1 0 1 0 2 Z0=120 TD=5n
SW1 0 1 3 0 inter
VCC 3 0 PULSE(0 5 0 1n 1n 500m)
VDD 4 0 DC 5
Rpullup 2 4 50k
D1 2 4 D1N4148
D2 0 2 D1N4148

.control
tran 10n 1u 0 1n
plot v(2)
.endc
.end
