Ouverture interrupteur sur ligne sans perte

.MODEL inter SW(RON=1m ROFF=10MEG VT=2.5 VH=.5)
SW1 0 1 3 0 inter
T1 1 0 2 0 Z0=120 TD=5n
VCC 3 0 PULSE(5 0 0 1n 1n 500m)
VDD 4 0 DC 5
Rpullup 2 4 50k

.control
tran 10n 1u 0 1n
plot v(2)
.endc
.end
