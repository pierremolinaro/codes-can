Ligne avec perte terminee par RC

.MODEL maLigne LTRA(R=70m L=600n C=41.7p G=0 LEN=1)
O1 0 1 0 2 maLigne
VCC 1 0 PULSE(0 5 0m 1n 1n 500m)
R1 0 2 120

.control
tran 10n 100n 0 1n
plot v(2)
.endc
.end
